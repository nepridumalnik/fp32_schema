`ifndef __CONST_SV__
`define __CONST_SV__

// Положительная бесконечность
`define P_INF32 32'h7F800000

// Ноль
`define ZERO32 32'h00000000

// Положительное не число
`define NAN32 32'h7FC00000

`endif
