typedef logic [31:0] Float32;
