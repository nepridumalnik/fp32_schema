`ifndef __TYPES_SV__
`define __TYPES_SV__

typedef logic [31:0] Float32;

`endif
